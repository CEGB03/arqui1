module Ej1( input logic x,
				output logic y);
		assign y = ~x;
endmodule 