module inversor(input logic x,
					output logic y);
	assign y= ~x;
endmodule