module Demo(input logic x,
				output logic y);
		assign y=~x;
endmodule 